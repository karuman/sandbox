module bot(bot_p1);
   input bot_p1;
   initial $monitor($stime ,, "bot_p1 = %b" , bot_p1);
endmodule
